
L1 N1P1 N1P2 0.1868u
E1_2 N1P3 N1P2 N2P1 N2P13 -0.3645
E1_3 N1P4 N1P3 N3P1 N3P13 -0.0311
E1_4 N1P5 N1P4 N4P1 N4P13 -0.0202
E1_5 N1P6 N1P5 N5P1 N5P13 -0.0121
E1_6 N1P7 N1P6 N6P1 N6P13 -0.0098
E1_7 N1P8 N1P7 N7P1 N7P13 -0.0015
E1_8 N1P9 N1P8 N8P1 N8P13 -0.0015
E1_9 N1P10 N1P9 N9P1 N9P13 -0.0024
E1_10 N1P11 N1P10 N10P1 N10P13 -0.0002
E1_11 N1P12 N1P11 N11P1 N11P13 -0.0687
E1_12 N1P13 N1P12 N12P1 N12P13 -0.3738
R1 N1P13 N2P1 R=1 LAPLACE=+1/{K1}/(-S*S/4/3.14^2)^0.25
.param K1=5.2884e-05
Ctt1_2 N1P1 N2P1 11.48p

L2 N2P1 N2P2 0.1490u
E2_1 N2P3 N2P2 N1P1 N1P13 -0.2909
E2_3 N2P4 N2P3 N3P1 N3P13 -0.3009
E2_4 N2P5 N2P4 N4P1 N4P13 -0.0189
E2_5 N2P6 N2P5 N5P1 N5P13 -0.0128
E2_6 N2P7 N2P6 N6P1 N6P13 -0.0094
E2_7 N2P8 N2P7 N7P1 N7P13 -0.0003
E2_8 N2P9 N2P8 N8P1 N8P13 0.0009
E2_9 N2P10 N2P9 N9P1 N9P13 0.0047
E2_10 N2P11 N2P10 N10P1 N10P13 -0.0527
E2_11 N2P12 N2P11 N11P1 N11P13 -0.2250
E2_12 N2P13 N2P12 N12P1 N12P13 -0.0548
R2 N2P13 N3P1 R=1 LAPLACE=+1/{K2}/(-S*S/4/3.14^2)^0.25
.param K2=4.9375e-05
Ctt2_3 N2P1 N3P1 10.69p

L3 N3P1 N3P2 0.1383u
E3_1 N3P3 N3P2 N1P1 N1P13 -0.0230
E3_2 N3P4 N3P3 N2P1 N2P13 -0.2793
E3_4 N3P5 N3P4 N4P1 N4P13 -0.3011
E3_5 N3P6 N3P5 N5P1 N5P13 -0.0188
E3_6 N3P7 N3P6 N6P1 N6P13 -0.0161
E3_7 N3P8 N3P7 N7P1 N7P13 -0.0006
E3_8 N3P9 N3P8 N8P1 N8P13 0.0049
E3_9 N3P10 N3P9 N9P1 N9P13 -0.0526
E3_10 N3P11 N3P10 N10P1 N10P13 -0.2244
E3_11 N3P12 N3P11 N11P1 N11P13 -0.0490
E3_12 N3P13 N3P12 N12P1 N12P13 -0.0001
R3 N3P13 N4P1 R=1 LAPLACE=+1/{K3}/(-S*S/4/3.14^2)^0.25
.param K3=4.5867e-05
Ctt3_4 N3P1 N4P1 9.90p

L4 N4P1 N4P2 0.1277u
E4_1 N4P3 N4P2 N1P1 N1P13 -0.0138
E4_2 N4P4 N4P3 N2P1 N2P13 -0.0162
E4_3 N4P5 N4P4 N3P1 N3P13 -0.2780
E4_5 N4P6 N4P5 N5P1 N5P13 -0.3021
E4_6 N4P7 N4P6 N6P1 N6P13 -0.0249
E4_7 N4P8 N4P7 N7P1 N7P13 0.0019
E4_8 N4P9 N4P8 N8P1 N8P13 -0.0527
E4_9 N4P10 N4P9 N9P1 N9P13 -0.2242
E4_10 N4P11 N4P10 N10P1 N10P13 -0.0485
E4_11 N4P12 N4P11 N11P1 N11P13 0.0040
E4_12 N4P13 N4P12 N12P1 N12P13 -0.0016
R4 N4P13 N5P1 R=1 LAPLACE=+1/{K4}/(-S*S/4/3.14^2)^0.25
.param K4=4.2358e-05
Ctt4_5 N4P1 N5P1 9.11p

L5 N5P1 N5P2 0.1172u
E5_1 N5P3 N5P2 N1P1 N1P13 -0.0076
E5_2 N5P4 N5P3 N2P1 N2P13 -0.0100
E5_3 N5P5 N5P4 N3P1 N3P13 -0.0159
E5_4 N5P6 N5P5 N4P1 N4P13 -0.2772
E5_6 N5P7 N5P6 N6P1 N6P13 -0.3125
E5_7 N5P8 N5P7 N7P1 N7P13 -0.0568
E5_8 N5P9 N5P8 N8P1 N8P13 -0.2243
E5_9 N5P10 N5P9 N9P1 N9P13 -0.0483
E5_10 N5P11 N5P10 N10P1 N10P13 0.0041
E5_11 N5P12 N5P11 N11P1 N11P13 0.0007
E5_12 N5P13 N5P12 N12P1 N12P13 -0.0009
R5 N5P13 N6P1 R=1 LAPLACE=+1/{K5}/(-S*S/4/3.14^2)^0.25
.param K5=3.8850e-05
Ctt5_6 N5P1 N6P1 8.33p

L6 N6P1 N6P2 0.1233u
E6_1 N6P3 N6P2 N1P1 N1P13 -0.0065
E6_2 N6P4 N6P3 N2P1 N2P13 -0.0078
E6_3 N6P5 N6P4 N3P1 N3P13 -0.0143
E6_4 N6P6 N6P5 N4P1 N4P13 -0.0240
E6_5 N6P7 N6P6 N5P1 N5P13 -0.3288
E6_7 N6P8 N6P7 N7P1 N7P13 -0.3573
E6_8 N6P9 N6P8 N8P1 N8P13 -0.0597
E6_9 N6P10 N6P9 N9P1 N9P13 0.0018
E6_10 N6P11 N6P10 N10P1 N10P13 -0.0006
E6_11 N6P12 N6P11 N11P1 N11P13 -0.0002
E6_12 N6P13 N6P12 N12P1 N12P13 -0.0010
R6 N6P13 N7P1 R=1 LAPLACE=+1/{K6}/(-S*S/4/3.14^2)^0.25
.param K6=3.5342e-05

L7 N7P1 N7P2 0.1233u
E7_1 N7P3 N7P2 N1P1 N1P13 -0.0010
E7_2 N7P4 N7P3 N2P1 N2P13 -0.0002
E7_3 N7P5 N7P4 N3P1 N3P13 -0.0006
E7_4 N7P6 N7P5 N4P1 N4P13 0.0018
E7_5 N7P7 N7P6 N5P1 N5P13 -0.0597
E7_6 N7P8 N7P7 N6P1 N6P13 -0.3573
E7_8 N7P9 N7P8 N8P1 N8P13 -0.3288
E7_9 N7P10 N7P9 N9P1 N9P13 -0.0240
E7_10 N7P11 N7P10 N10P1 N10P13 -0.0143
E7_11 N7P12 N7P11 N11P1 N11P13 -0.0078
E7_12 N7P13 N7P12 N12P1 N12P13 -0.0065
R7 N7P13 N8P1 R=1 LAPLACE=+1/{K7}/(-S*S/4/3.14^2)^0.25
.param K7=3.5342e-05
Ctt7_8 N7P1 N8P1 8.33p

L8 N8P1 N8P2 0.1172u
E8_1 N8P3 N8P2 N1P1 N1P13 -0.0009
E8_2 N8P4 N8P3 N2P1 N2P13 0.0007
E8_3 N8P5 N8P4 N3P1 N3P13 0.0041
E8_4 N8P6 N8P5 N4P1 N4P13 -0.0483
E8_5 N8P7 N8P6 N5P1 N5P13 -0.2243
E8_6 N8P8 N8P7 N6P1 N6P13 -0.0568
E8_7 N8P9 N8P8 N7P1 N7P13 -0.3125
E8_9 N8P10 N8P9 N9P1 N9P13 -0.2772
E8_10 N8P11 N8P10 N10P1 N10P13 -0.0159
E8_11 N8P12 N8P11 N11P1 N11P13 -0.0100
E8_12 N8P13 N8P12 N12P1 N12P13 -0.0076
R8 N8P13 N9P1 R=1 LAPLACE=+1/{K8}/(-S*S/4/3.14^2)^0.25
.param K8=3.8850e-05
Ctt8_9 N8P1 N9P1 9.11p

L9 N9P1 N9P2 0.1277u
E9_1 N9P3 N9P2 N1P1 N1P13 -0.0016
E9_2 N9P4 N9P3 N2P1 N2P13 0.0040
E9_3 N9P5 N9P4 N3P1 N3P13 -0.0485
E9_4 N9P6 N9P5 N4P1 N4P13 -0.2242
E9_5 N9P7 N9P6 N5P1 N5P13 -0.0527
E9_6 N9P8 N9P7 N6P1 N6P13 0.0019
E9_7 N9P9 N9P8 N7P1 N7P13 -0.0249
E9_8 N9P10 N9P9 N8P1 N8P13 -0.3021
E9_10 N9P11 N9P10 N10P1 N10P13 -0.2780
E9_11 N9P12 N9P11 N11P1 N11P13 -0.0162
E9_12 N9P13 N9P12 N12P1 N12P13 -0.0138
R9 N9P13 N10P1 R=1 LAPLACE=+1/{K9}/(-S*S/4/3.14^2)^0.25
.param K9=4.2358e-05
Ctt9_10 N9P1 N10P1 9.90p

L10 N10P1 N10P2 0.1383u
E10_1 N10P3 N10P2 N1P1 N1P13 -0.0001
E10_2 N10P4 N10P3 N2P1 N2P13 -0.0490
E10_3 N10P5 N10P4 N3P1 N3P13 -0.2244
E10_4 N10P6 N10P5 N4P1 N4P13 -0.0526
E10_5 N10P7 N10P6 N5P1 N5P13 0.0049
E10_6 N10P8 N10P7 N6P1 N6P13 -0.0006
E10_7 N10P9 N10P8 N7P1 N7P13 -0.0161
E10_8 N10P10 N10P9 N8P1 N8P13 -0.0188
E10_9 N10P11 N10P10 N9P1 N9P13 -0.3011
E10_11 N10P12 N10P11 N11P1 N11P13 -0.2793
E10_12 N10P13 N10P12 N12P1 N12P13 -0.0230
R10 N10P13 N11P1 R=1 LAPLACE=+1/{K10}/(-S*S/4/3.14^2)^0.25
.param K10=4.5867e-05
Ctt10_11 N10P1 N11P1 10.69p

L11 N11P1 N11P2 0.1490u
E11_1 N11P3 N11P2 N1P1 N1P13 -0.0548
E11_2 N11P4 N11P3 N2P1 N2P13 -0.2250
E11_3 N11P5 N11P4 N3P1 N3P13 -0.0527
E11_4 N11P6 N11P5 N4P1 N4P13 0.0047
E11_5 N11P7 N11P6 N5P1 N5P13 0.0009
E11_6 N11P8 N11P7 N6P1 N6P13 -0.0003
E11_7 N11P9 N11P8 N7P1 N7P13 -0.0094
E11_8 N11P10 N11P9 N8P1 N8P13 -0.0128
E11_9 N11P11 N11P10 N9P1 N9P13 -0.0189
E11_10 N11P12 N11P11 N10P1 N10P13 -0.3009
E11_12 N11P13 N11P12 N12P1 N12P13 -0.2909
R11 N11P13 N12P1 R=1 LAPLACE=+1/{K11}/(-S*S/4/3.14^2)^0.25
.param K11=4.9375e-05
Ctt11_12 N11P1 N12P1 11.48p

L12 N12P1 N12P2 0.1868u
E12_1 N12P3 N12P2 N1P1 N1P13 -0.3738
E12_2 N12P4 N12P3 N2P1 N2P13 -0.0687
E12_3 N12P5 N12P4 N3P1 N3P13 -0.0002
E12_4 N12P6 N12P5 N4P1 N4P13 -0.0024
E12_5 N12P7 N12P6 N5P1 N5P13 -0.0015
E12_6 N12P8 N12P7 N6P1 N6P13 -0.0015
E12_7 N12P9 N12P8 N7P1 N7P13 -0.0098
E12_8 N12P10 N12P9 N8P1 N8P13 -0.0121
E12_9 N12P11 N12P10 N9P1 N9P13 -0.0202
E12_10 N12P12 N12P11 N10P1 N10P13 -0.0311
E12_11 N12P13 N12P12 N11P1 N11P13 -0.3645
R12 N12P13 N13P1 R=1 LAPLACE=+1/{K12}/(-S*S/4/3.14^2)^0.25
.param K12=5.2884e-05

Cdd1_12 N1P1 N12P1 11.87p
Cdd2_11 N2P1 N11P1 11.08p
Cdd3_10 N3P1 N10P1 10.30p
Cdd4_9 N4P1 N9P1 9.51p
Cdd5_8 N5P1 N8P1 8.72p
Cdd6_7 N6P1 N7P1 7.93p

V1 In 0 AC 10
Rin In N1P1 50
Rout N13P1 0 50
.print V(N13P1)
.print V(In)

.ac dec 1000 10 200000k
.backanno
.end
